module tb_linx_cpu_pyc;
  logic clk;
  logic rst;

  logic [63:0] boot_pc = 64'h0000_0000_0001_0000;
  logic [63:0] boot_sp = 64'h0000_0000_0002_0000;

  logic halted;
  logic [63:0] pc;
  logic [2:0] stage;
  logic [63:0] cycles;
  logic [63:0] a0;
  logic [63:0] a1;
  logic [63:0] ra;
  logic [63:0] sp;
  logic [2:0] br_kind;
  logic [63:0] if_window;
  logic [11:0] wb_op;
  logic [5:0] wb_regdst;
  logic [63:0] wb_value;
  logic commit_cond;
  logic [63:0] commit_tgt;

  logic [31:0] exit_code;
  logic uart_valid;
  logic [7:0] uart_byte;
  logic irq;
  logic [63:0] irq_vector;

  // Pipeview (Konata) stage hooks (exported as optional debug ports).
  logic if0_valid;
  logic [63:0] if0_pc;
  logic if1_valid;
  logic [63:0] if1_pc;
  logic ifid0_valid;
  logic [63:0] ifid0_pc;
  logic ifid1_valid;
  logic [63:0] ifid1_pc;
  logic idex0_valid;
  logic [63:0] idex0_pc;
  logic idex1_valid;
  logic [63:0] idex1_pc;
  logic exmem0_valid;
  logic [63:0] exmem0_pc;
  logic exmem1_valid;
  logic [63:0] exmem1_pc;
  logic wb0_valid;
  logic wb1_valid;
  logic [63:0] wb0_pc;
  logic [63:0] wb1_pc;
  logic [11:0] wb0_op;
  logic [11:0] wb1_op;

  // Generated by pyc-compile: module linx_cpu_pyc
  linx_cpu_pyc dut (
      .clk(clk),
      .rst(rst),
      .boot_pc(boot_pc),
      .boot_sp(boot_sp),
      .irq(irq),
      .irq_vector(irq_vector),
      .host_wvalid(1'b0),
      .host_waddr(64'd0),
      .host_wdata(64'd0),
      .host_wstrb(8'd0),
      .halted(halted),
      .exit_code(exit_code),
      .uart_valid(uart_valid),
      .uart_byte(uart_byte),
      .pc(pc),
      .stage(stage),
      .cycles(cycles),
      .a0(a0),
      .a1(a1),
      .ra(ra),
      .sp(sp),
      .br_kind(br_kind),
      .if_window(if_window),
      .if0_valid(if0_valid),
      .if0_pc(if0_pc),
      .if1_valid(if1_valid),
      .if1_pc(if1_pc),
      .ifid0_valid(ifid0_valid),
      .ifid0_pc(ifid0_pc),
      .ifid1_valid(ifid1_valid),
      .ifid1_pc(ifid1_pc),
      .idex0_valid(idex0_valid),
      .idex0_pc(idex0_pc),
      .idex1_valid(idex1_valid),
      .idex1_pc(idex1_pc),
      .exmem0_valid(exmem0_valid),
      .exmem0_pc(exmem0_pc),
      .exmem1_valid(exmem1_valid),
      .exmem1_pc(exmem1_pc),
      .wb0_valid(wb0_valid),
      .wb0_pc(wb0_pc),
      .wb0_op(wb0_op),
      .wb1_valid(wb1_valid),
      .wb1_pc(wb1_pc),
      .wb1_op(wb1_op),
      .wb_op(wb_op),
      .wb_regdst(wb_regdst),
      .wb_value(wb_value),
      .commit_cond(commit_cond),
      .commit_tgt(commit_tgt)
  );

  always #5 clk = ~clk;

  function automatic logic [31:0] mem_read32(input int unsigned addr);
    mem_read32 = {dut.dmem.mem[addr + 3], dut.dmem.mem[addr + 2], dut.dmem.mem[addr + 1], dut.dmem.mem[addr + 0]};
  endfunction

  string memh_path;
  int unsigned expected;
  int unsigned expected_exit;
  bit do_memcheck;
  string vcd_path;
  string log_path;
  int log_fd;
  bit log_cycles;
  string konata_path;
  int konata_fd;
  bit konata_on;
  longint unsigned konata_cur_cycle;
  longint unsigned konata_next_id;
  typedef struct {
    bit v;
    longint unsigned id;
    longint unsigned pc;
  } slot_t;
  slot_t prev_if[2];
  slot_t prev_id[2];
  slot_t prev_ex[2];
  slot_t prev_mem[2];
  slot_t prev_wb[2];
  slot_t cur_if[2];
  slot_t cur_id[2];
  slot_t cur_ex[2];
  slot_t cur_mem[2];
  slot_t cur_wb[2];
  int i;
  logic [31:0] got;

  task automatic konata_at_cycle(input longint unsigned cyc);
    if (!konata_on)
      return;
    if (cyc < konata_cur_cycle)
      return;
    if (cyc == konata_cur_cycle)
      return;
    $fdisplay(konata_fd, "C\t%0d", (cyc - konata_cur_cycle));
    konata_cur_cycle = cyc;
  endtask

  task automatic konata_insn(input longint unsigned file_id, input longint unsigned sim_id, input longint unsigned thread_id);
    if (konata_on)
      $fdisplay(konata_fd, "I\t%0d\t%0d\t%0d", file_id, sim_id, thread_id);
  endtask

  task automatic konata_label(input longint unsigned id, input int kind, input string msg);
    if (konata_on)
      $fdisplay(konata_fd, "L\t%0d\t%0d\t%s", id, kind, msg);
  endtask

  task automatic konata_stage_start(input longint unsigned id, input int lane, input string stage);
    if (konata_on)
      $fdisplay(konata_fd, "S\t%0d\t%0d\t%s", id, lane, stage);
  endtask

  task automatic konata_stage_end(input longint unsigned id, input int lane, input string stage);
    if (konata_on)
      $fdisplay(konata_fd, "E\t%0d\t%0d\t%s", id, lane, stage);
  endtask

  task automatic konata_retire(input longint unsigned id, input longint unsigned retire_id, input int kind);
    if (konata_on)
      $fdisplay(konata_fd, "R\t%0d\t%0d\t%0d", id, retire_id, kind);
  endtask

  task automatic pv_alloc_id(input longint unsigned pc, input int lane, output longint unsigned id);
    id = konata_next_id;
    konata_next_id++;
    konata_insn(id, pc, 0);
    konata_label(id, 0, $sformatf("pc=0x%016x lane=%0d", pc, lane));
  endtask

  task automatic pv_assign_slot(
      input bit valid,
      input longint unsigned pc,
      input slot_t prev_same,
      input slot_t prev_from,
      input bit allow_from,
      input int lane,
      output slot_t out);
    out.v = valid;
    out.pc = pc;
    out.id = 0;
    if (!valid)
      return;
    if (prev_same.v && prev_same.pc == pc) begin
      out.id = prev_same.id;
      return;
    end
    if (allow_from && prev_from.v && prev_from.pc == pc) begin
      out.id = prev_from.id;
      return;
    end
    pv_alloc_id(pc, lane, out.id);
  endtask

  task automatic pv_stage_update(input slot_t prev_s, input slot_t cur_s, input int lane, input string stage, input bit retire_on_end);
    if (!konata_on)
      return;
    if (prev_s.v && (!cur_s.v || (cur_s.id != prev_s.id))) begin
      konata_stage_end(prev_s.id, lane, stage);
      if (retire_on_end)
        konata_retire(prev_s.id, prev_s.id, 0);
    end
    if (cur_s.v && (!prev_s.v || (cur_s.id != prev_s.id))) begin
      konata_stage_start(cur_s.id, lane, stage);
    end
  endtask

  initial begin
    clk = 1'b0;
    rst = 1'b1;
    irq = 1'b0;
    irq_vector = 64'd0;
    if (!$value$plusargs("memh=%s", memh_path)) begin
      memh_path = "designs/examples/linx_cpu/programs/test_or.memh";
    end
    if (!$value$plusargs("expected=%h", expected)) begin
      expected = 32'h0000_ff00;
    end
    if (!$value$plusargs("expected_exit=%h", expected_exit)) begin
      expected_exit = 32'h0000_0000;
    end
    do_memcheck = !$test$plusargs("no_memcheck");

    // Tracing / logging (default: enabled; disable with +notrace / +nolog).
    vcd_path = ".pycircuit_out/examples/linx_cpu_pyc/tb_linx_cpu_pyc_sv.vcd";
    log_path = ".pycircuit_out/examples/linx_cpu_pyc/tb_linx_cpu_pyc_sv.log";
    konata_path = ".pycircuit_out/examples/linx_cpu_pyc/tb_linx_cpu_pyc_sv.konata";
    void'($value$plusargs("vcd=%s", vcd_path));
    void'($value$plusargs("log=%s", log_path));
    void'($value$plusargs("konata=%s", konata_path));
    log_cycles = $test$plusargs("logcycles");
    konata_on = !$test$plusargs("nokonata");
    konata_fd = 0;
    konata_next_id = 1;
    if (konata_on) begin
      konata_fd = $fopen(konata_path, "w");
      if (konata_fd == 0) begin
        $display("WARN: failed to open Konata log: %s", konata_path);
        konata_on = 0;
      end
    end

    if (!$test$plusargs("notrace")) begin
      $display("tb_linx_cpu_pyc: dumping VCD to %s", vcd_path);
      $dumpfile(vcd_path);
      $dumpvars(0, tb_linx_cpu_pyc);
    end

    if (!$test$plusargs("nolog")) begin
      log_fd = $fopen(log_path, "w");
      $fdisplay(log_fd, "tb_linx_cpu_pyc(SV): memh=%s expected=0x%08x", memh_path, expected);
      $fdisplay(log_fd, "cycle,time,halted,stage,pc,cycles");
    end else begin
      log_fd = 0;
    end

    $display("tb_linx_cpu_pyc: memh=%s expected=0x%08x expected_exit=0x%08x", memh_path, expected, expected_exit);

    // Bring-up model has separate I$ + D$ byte memories. Load the image into both.
    $readmemh(memh_path, dut.imem.mem);
    $readmemh(memh_path, dut.dmem.mem);

    repeat (5) @(posedge clk);
    rst = 1'b0;

    if (konata_on) begin
      $fdisplay(konata_fd, "Kanata\t0004");
      $fdisplay(konata_fd, "C=\t%0d", cycles);
      konata_cur_cycle = cycles;
      for (int lane = 0; lane < 2; lane++) begin
        prev_if[lane].v = 0;
        prev_if[lane].id = 0;
        prev_if[lane].pc = 0;
        prev_id[lane].v = 0;
        prev_id[lane].id = 0;
        prev_id[lane].pc = 0;
        prev_ex[lane].v = 0;
        prev_ex[lane].id = 0;
        prev_ex[lane].pc = 0;
        prev_mem[lane].v = 0;
        prev_mem[lane].id = 0;
        prev_mem[lane].pc = 0;
        prev_wb[lane].v = 0;
        prev_wb[lane].id = 0;
        prev_wb[lane].pc = 0;
      end
    end

    i = 0;
    while (i < 200000 && !halted) begin
      @(posedge clk);
      if (konata_on) begin
        konata_at_cycle(cycles);

        // Lane 0.
        pv_assign_slot(if0_valid, if0_pc, prev_if[0], prev_if[0], 0, 0, cur_if[0]);
        pv_assign_slot(ifid0_valid, ifid0_pc, prev_id[0], prev_if[0], 1, 0, cur_id[0]);
        pv_assign_slot(idex0_valid, idex0_pc, prev_ex[0], prev_id[0], 1, 0, cur_ex[0]);
        pv_assign_slot(exmem0_valid, exmem0_pc, prev_mem[0], prev_ex[0], 1, 0, cur_mem[0]);
        pv_assign_slot(wb0_valid, wb0_pc, prev_wb[0], prev_mem[0], 1, 0, cur_wb[0]);

        pv_stage_update(prev_if[0], cur_if[0], 0, "IF", 0);
        pv_stage_update(prev_id[0], cur_id[0], 0, "ID", 0);
        pv_stage_update(prev_ex[0], cur_ex[0], 0, "EX", 0);
        pv_stage_update(prev_mem[0], cur_mem[0], 0, "MEM", 0);
        pv_stage_update(prev_wb[0], cur_wb[0], 0, "WB", 1);
        if (cur_wb[0].v && (!prev_wb[0].v || (cur_wb[0].id != prev_wb[0].id)))
          konata_label(cur_wb[0].id, 1, $sformatf("wb op=%0d", wb0_op));

        prev_if[0] = cur_if[0];
        prev_id[0] = cur_id[0];
        prev_ex[0] = cur_ex[0];
        prev_mem[0] = cur_mem[0];
        prev_wb[0] = cur_wb[0];

        // Lane 1.
        pv_assign_slot(if1_valid, if1_pc, prev_if[1], prev_if[1], 0, 1, cur_if[1]);
        pv_assign_slot(ifid1_valid, ifid1_pc, prev_id[1], prev_if[1], 1, 1, cur_id[1]);
        pv_assign_slot(idex1_valid, idex1_pc, prev_ex[1], prev_id[1], 1, 1, cur_ex[1]);
        pv_assign_slot(exmem1_valid, exmem1_pc, prev_mem[1], prev_ex[1], 1, 1, cur_mem[1]);
        pv_assign_slot(wb1_valid, wb1_pc, prev_wb[1], prev_mem[1], 1, 1, cur_wb[1]);

        pv_stage_update(prev_if[1], cur_if[1], 1, "IF", 0);
        pv_stage_update(prev_id[1], cur_id[1], 1, "ID", 0);
        pv_stage_update(prev_ex[1], cur_ex[1], 1, "EX", 0);
        pv_stage_update(prev_mem[1], cur_mem[1], 1, "MEM", 0);
        pv_stage_update(prev_wb[1], cur_wb[1], 1, "WB", 1);
        if (cur_wb[1].v && (!prev_wb[1].v || (cur_wb[1].id != prev_wb[1].id)))
          konata_label(cur_wb[1].id, 1, $sformatf("wb op=%0d", wb1_op));

        prev_if[1] = cur_if[1];
        prev_id[1] = cur_id[1];
        prev_ex[1] = cur_ex[1];
        prev_mem[1] = cur_mem[1];
        prev_wb[1] = cur_wb[1];
      end
      if (uart_valid) begin
        $write("%c", uart_byte);
      end
      if (log_fd != 0 && log_cycles) begin
        $fdisplay(log_fd, "%0d,%0t,%0b,%0d,0x%016x,%0d", i, $time, halted, stage, pc, cycles);
      end
      i++;
    end

    if (!halted) begin
      $fatal(1, "FAIL: did not halt (pc=0x%016x cycles=%0d)", pc, cycles);
    end

    if (exit_code !== expected_exit[31:0]) begin
      $fatal(1, "FAIL: exit_code=0x%08x expected_exit=0x%08x", exit_code, expected_exit[31:0]);
    end

    got = mem_read32(32'h0000_0100);
    if (do_memcheck && got !== expected[31:0]) begin
      $fatal(1, "FAIL: mem[0x100]=0x%08x expected=0x%08x", got, expected[31:0]);
    end

    if (log_fd != 0) begin
      $fdisplay(log_fd, "PASS: mem[0x100]=0x%08x cycles=%0d pc=0x%016x", got, cycles, pc);
      $fclose(log_fd);
    end

    if (konata_fd != 0) begin
      $fclose(konata_fd);
    end

    $display("PASS: mem[0x100]=0x%08x cycles=%0d", got, cycles);
    $finish;
  end

endmodule
